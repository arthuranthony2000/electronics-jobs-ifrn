CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
10 0 1 90 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
48 C:\Program Files\CircuitMaker 2000 Trial\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
35
7 Ground~
168 1032 89 0 1 3
0 2
0
0 0 53360 180
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9274 0 0
2
5.89786e-315 0
0
2 +V
167 1232 49 0 1 3
0 13
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V9
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4197 0 0
2
5.89786e-315 0
0
9 CA 7-Seg~
184 1232 93 0 18 19
10 12 11 10 9 8 7 6 33 13
0 0 2 0 0 2 0 2 1
0
0 0 21088 0
6 BLUECA
13 -41 55 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
7363 0 0
2
5.89786e-315 0
0
6 74LS47
187 1097 180 0 14 29
0 2 3 4 5 34 35 6 7 8
9 10 11 12 36
0
0 0 4848 0
6 74LS47
-21 -60 21 -52
2 U6
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
4319 0 0
2
5.89786e-315 0
0
7 Pulser~
4 1004 565 0 10 12
0 37 38 14 39 0 0 10 10 6
8
0
0 0 4656 180
0
2 V8
-7 -29 7 -21
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3919 0 0
2
42762.9 0
0
9 2-In AND~
219 674 250 0 3 22
0 17 4 16
0
0 0 624 90
6 74LS08
-21 -24 21 -16
3 U5A
16 -5 37 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
7852 0 0
2
42762.9 1
0
8 2-In OR~
219 389 406 0 3 22
0 21 20 19
0
0 0 624 180
6 74LS32
-21 -24 21 -16
3 U3C
1 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
9310 0 0
2
42762.9 2
0
9 2-In AND~
219 466 430 0 3 22
0 5 18 21
0
0 0 624 180
6 74LS08
-21 -24 21 -16
3 U4D
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
8989 0 0
2
42762.9 3
0
9 2-In AND~
219 461 380 0 3 22
0 17 3 20
0
0 0 624 180
6 74LS08
-21 -24 21 -16
3 U4C
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
3598 0 0
2
42762.9 4
0
2 +V
167 447 190 0 1 3
0 22
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V7
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3842 0 0
2
42762.9 5
0
8 2-In OR~
219 202 340 0 3 22
0 15 3 23
0
0 0 624 180
6 74LS32
-21 -24 21 -16
3 U3B
1 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
7145 0 0
2
42762.9 6
0
7 Ground~
168 801 482 0 1 3
0 2
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6598 0 0
2
42762.9 7
0
7 Ground~
168 483 483 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9435 0 0
2
42762.9 8
0
7 Ground~
168 209 492 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3397 0 0
2
42762.9 9
0
4 LED~
171 901 455 0 2 2
10 18 2
0
0 0 864 0
4 LED0
17 0 45 8
2 D6
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
5438 0 0
2
42762.9 10
0
4 LED~
171 577 455 0 2 2
10 15 2
0
0 0 864 0
4 LED0
17 0 45 8
2 D5
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3222 0 0
2
42762.9 11
0
4 LED~
171 297 451 0 2 2
10 17 2
0
0 0 864 0
4 LED0
17 0 45 8
2 D4
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3733 0 0
2
42762.9 12
0
9 2-In AND~
219 182 60 0 3 22
0 15 3 24
0
0 0 624 180
6 74LS08
-21 -24 21 -16
3 U4B
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
3856 0 0
2
42762.9 13
0
9 2-In AND~
219 189 112 0 3 22
0 4 18 25
0
0 0 624 180
6 74LS08
-21 -24 21 -16
3 U4A
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
5122 0 0
2
42762.9 14
0
8 2-In OR~
219 112 88 0 3 22
0 25 24 26
0
0 0 624 180
6 74LS32
-21 -24 21 -16
3 U3A
1 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3597 0 0
2
42762.9 15
0
2 +V
167 775 276 0 1 3
0 27
0
0 0 54256 180
3 10V
6 -2 27 6
2 V6
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6559 0 0
2
42762.9 16
0
2 +V
167 775 179 0 1 3
0 28
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7392 0 0
2
42762.9 17
0
2 +V
167 497 271 0 1 3
0 29
0
0 0 54256 180
3 10V
6 -2 27 6
2 V4
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4519 0 0
2
42762.9 18
0
2 +V
167 497 174 0 1 3
0 30
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3878 0 0
2
42762.9 19
0
2 +V
167 240 272 0 1 3
0 32
0
0 0 54256 180
3 10V
6 -2 27 6
2 V2
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6230 0 0
2
42762.9 20
0
2 +V
167 240 175 0 1 3
0 31
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5407 0 0
2
42762.9 21
0
7 Ground~
168 814 26 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9885 0 0
2
42762.9 22
0
7 Ground~
168 490 28 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5899 0 0
2
42762.9 23
0
7 Ground~
168 232 30 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7294 0 0
2
42762.9 24
0
4 LED~
171 897 28 0 2 2
10 3 2
0
0 0 864 180
4 LED0
16 0 44 8
2 D3
23 -10 37 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
5851 0 0
2
42762.9 25
0
4 LED~
171 577 29 0 2 2
10 4 2
0
0 0 864 180
4 LED0
16 0 44 8
2 D2
23 -10 37 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
6635 0 0
2
42762.9 26
0
4 LED~
171 307 31 0 2 2
10 5 2
0
0 0 864 180
4 LED0
16 0 44 8
2 D1
23 -10 37 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3726 0 0
2
42762.9 27
0
6 74112~
219 775 250 0 7 32
0 28 16 14 15 27 18 3
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 1 2 0
1 U
317 0 0
2
42762.9 28
0
6 74112~
219 497 245 0 7 32
0 30 22 14 19 29 15 4
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U1B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 2 1 0
1 U
5827 0 0
2
42762.9 29
0
6 74112~
219 240 246 0 7 32
0 31 26 14 23 32 17 5
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U1A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 1 1 0
1 U
7681 0 0
2
42762.9 30
0
55
2 0 3 0 0 8192 0 4 0 0 53 3
1065 153
1065 158
899 158
3 0 4 0 0 4224 0 4 0 0 54 2
1065 162
579 162
4 0 5 0 0 12416 0 4 0 0 55 4
1065 171
782 171
782 157
309 157
1 1 2 0 0 8192 0 4 1 0 0 3
1065 144
1032 144
1032 97
7 7 6 0 0 4224 0 4 3 0 0 3
1135 144
1247 144
1247 129
8 6 7 0 0 4224 0 4 3 0 0 3
1135 153
1241 153
1241 129
9 5 8 0 0 4224 0 4 3 0 0 3
1135 162
1235 162
1235 129
10 4 9 0 0 4224 0 4 3 0 0 3
1135 171
1229 171
1229 129
11 3 10 0 0 4224 0 4 3 0 0 3
1135 180
1223 180
1223 129
12 2 11 0 0 4224 0 4 3 0 0 3
1135 189
1217 189
1217 129
13 1 12 0 0 4224 0 4 3 0 0 3
1135 198
1211 198
1211 129
1 9 13 0 0 4224 0 2 3 0 0 2
1232 58
1232 57
3 0 14 0 0 8192 0 33 0 0 15 3
745 223
742 223
742 572
3 0 14 0 0 0 0 34 0 0 15 7
467 218
463 218
463 361
486 361
486 411
436 411
436 572
3 3 14 0 0 12416 0 35 5 0 0 4
210 219
100 219
100 572
980 572
4 0 15 0 0 8192 0 33 0 0 39 4
751 232
723 232
723 397
577 397
3 2 16 0 0 8320 0 6 33 0 0 3
673 226
673 214
751 214
2 0 4 0 0 0 0 6 0 0 54 5
682 271
682 299
593 299
593 177
579 177
1 0 17 0 0 8320 0 6 0 0 40 3
664 271
664 279
297 279
2 0 3 0 0 4096 0 9 0 0 53 4
479 371
851 371
851 171
899 171
1 0 17 0 0 0 0 9 0 0 40 4
479 389
532 389
532 290
297 290
2 0 18 0 0 4096 0 8 0 0 38 2
484 421
901 421
1 0 5 0 0 0 0 8 0 0 55 6
484 439
505 439
505 308
386 308
386 170
309 170
3 4 19 0 0 8320 0 7 34 0 0 4
362 406
354 406
354 227
473 227
2 3 20 0 0 8320 0 7 9 0 0 4
408 397
424 397
424 380
434 380
1 3 21 0 0 4224 0 7 8 0 0 4
408 415
424 415
424 430
439 430
1 2 22 0 0 8320 0 10 34 0 0 3
447 199
447 209
473 209
2 0 3 0 0 4096 0 11 0 0 53 4
221 331
873 331
873 151
899 151
1 0 15 0 0 4096 0 11 0 0 39 2
221 349
577 349
3 4 23 0 0 8320 0 11 35 0 0 4
175 340
168 340
168 228
216 228
2 0 3 0 0 4224 0 18 0 0 53 2
200 51
899 51
1 0 15 0 0 4224 0 18 0 0 39 4
200 69
610 69
610 319
577 319
2 0 18 0 0 4224 0 19 0 0 38 4
207 103
934 103
934 372
901 372
1 0 4 0 0 0 0 19 0 0 54 2
207 121
579 121
1 2 2 0 0 8320 0 12 15 0 0 4
801 476
801 471
901 471
901 465
1 2 2 0 0 0 0 13 16 0 0 4
483 477
483 473
577 473
577 465
1 2 2 0 0 0 0 14 17 0 0 4
209 486
209 469
297 469
297 461
6 1 18 0 0 0 0 33 15 0 0 3
805 232
901 232
901 445
6 1 15 0 0 0 0 34 16 0 0 3
527 227
577 227
577 445
6 1 17 0 0 0 0 35 17 0 0 3
270 228
297 228
297 441
2 3 24 0 0 4224 0 20 18 0 0 4
131 79
154 79
154 60
155 60
1 3 25 0 0 4224 0 20 19 0 0 4
131 97
156 97
156 112
162 112
3 2 26 0 0 12416 0 20 35 0 0 4
85 88
80 88
80 210
216 210
1 5 27 0 0 4224 0 21 33 0 0 2
775 261
775 262
1 1 28 0 0 4224 0 22 33 0 0 2
775 188
775 187
1 5 29 0 0 4224 0 23 34 0 0 2
497 256
497 257
1 1 30 0 0 4224 0 24 34 0 0 2
497 183
497 182
1 1 31 0 0 4224 0 26 35 0 0 2
240 184
240 183
1 5 32 0 0 4224 0 25 35 0 0 2
240 257
240 258
1 2 2 0 0 0 0 27 30 0 0 4
814 20
814 10
899 10
899 18
1 2 2 0 0 0 0 29 32 0 0 4
232 24
232 13
309 13
309 21
1 2 2 0 0 0 0 28 31 0 0 4
490 22
490 11
579 11
579 19
7 1 3 0 0 0 0 33 30 0 0 3
799 214
899 214
899 38
7 1 4 0 0 0 0 34 31 0 0 3
521 209
579 209
579 39
7 1 5 0 0 0 0 35 32 0 0 3
264 210
309 210
309 41
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
